package switch_pkg; 
//	`include "env_config.sv"
//	`include "

	
	import uvm_pkg::*;
	`include "uvm_macros.svh"
`include "src_trans.sv"
//`include "ram_wr_agent_config.sv"
//`include "ram_rd_agent_config.sv"
`include "env_config.sv"
`include "src_driver.sv"
`include "src_monitor.sv"
`include "src_sequencer.sv"
`include "src_agent.sv"
`include "src_seq.sv"

`include "dest_trans.sv"
`include "dest_monitor.sv"
//`include "dest_sequencer.sv"
//`include "ram_rd_seqs.sv"
//`include "ram_rd_driver.sv"
`include "dest_agent.sv"
//`include "ram_rd_agt_top.sv"

//`include "ram_virtual_sequencer.sv"
//`include "ram_virtual_seqs.sv"
//`include "ram_scoreboard.sv"

`include "environment.sv"


`include "test.sv"
endpackage
